library ieee;

entity contador4 is
port (
clock: in bit ;
zera : in bit ;
conta : in bit ;
Q : out bit_vector ( 3 downto 0 ) ;
fim : out bit
) ;
end entity contador4 ;

architecture counter of contador4 is
    signal 

    if zera == 1 then
        Q <= "0000";
    else if 
        Q <= bit_vector(Q + '1') ;
begin

end architecture;